netcdf hru_attri {
dimensions:
	hru_id = 5 ;
	gru_id = 1 ;

variables:

data:


group: gru {
dimensions:
	gru_id = 1 ;

variables:
	int gru_id(gru_id) ;
		gru_id:long_name = "index of group of response unit (GRU)" ;
	int gru_start_id(gru_id) ;
		gru_start_id:long_name = "the index (hru_id) for the first hru in a gru " ;
	int gru_hCount(gru_id) ;
		gru_hCount:long_name = "the total number of hrus in a gru" ;

// group attributes:
	  :data_provider = "/home/huanwu/summa/fork/summa/setup_tools/input/" ;
	  :data_reference = "/home/huanwu/summa/fork/summa/setup_tools/output/" ;
data:

 gru_id = 1 ;

 gru_start_id = 1 ;

 gru_hCount = 5 ;

}

group: local_types {
dimensions:
	hru_id = 5 ;

variables:
	int hru_id(hru_id) ;
		hru_id:long_name = "index of hydrological response units (HRU)" ;
  	int vegTypeIndex(hru_id) ;
  		vegTypeIndex:long_name = "index defining vegetation type" ;
  		vegTypeIndex:units = "-" ;
  	int soilTypeIndex(hru_id) ;
  		soilTypeIndex:long_name = "index defining soil type" ;
  		soilTypeIndex:units = "-" ;
  	int slopeTypeIndex(hru_id) ;
  		slopeTypeIndex:long_name = "index defining slope" ;
  		slopeTypeIndex:units = "-" ;
  	int downHRUindex(hru_id) ;
  		downHRUindex:long_name = "index of downslope HRU (0 = basin outlet)" ;
  		downHRUindex:units = "-" ;
  	int GRUindex(hru_id) ;
  		GRUindex:long_name = "index of GRU to which the HRU belongs" ;
  		GRUindex:units = "-" ;

// group attributes:
	  :data_provider = "/home/huanwu/summa/fork/summa/setup_tools/input/" ;
	  :data_reference = "/home/huanwu/summa/fork/summa/setup_tools/output/" ;
data:

   hru_id = 1, 2, 3, 4, 5 ;

   vegTypeIndex = 11, 11, 11, 11, 11 ;

   soilTypeIndex = 8, 8, 8, 8, 8 ;

   slopeTypeIndex = 1, 1, 1, 1, 1 ;

   downHRUindex = 0, 0, 0, 0, 0 ;

   GRUindex = 1, 1, 1, 1, 1 ;

}

group: hru_attributes {
  dimensions:
  	hru_id = 5 ;
  variables:
  	double HRUarea(hru_id) ;
  		HRUarea:long_name = "area of each HRU" ;
  		HRUarea:units = "m^2" ;
  	double latitude(hru_id) ;
  		latitude:long_name = "latitude of HRU\'s centriod point" ;
  		latitude:units = "decimal degree north" ;
  	double longitude(hru_id) ;
  		longitude:long_name = "longitude of HRU\'s centriod point" ;
  		longitude:units = "decimal degree east" ;
  	double elevation(hru_id) ;
  		elevation:long_name = "elevation of HRU\'s centriod point" ;
  		elevation:units = "m" ;
  	double tan_slope(hru_id) ;
  		tan_slope:long_name = "average tangent slope of HRU" ;
  		tan_slope:units = "m m-1" ;
  	double contourLength(hru_id) ;
  		contourLength:long_name = "contourLength of HRU" ;
  		contourLength:units = "m" ;
  	double mHeight(hru_id) ;
  		mHeight:long_name = "measurement height above bare ground" ;
  		mHeight:units = "m" ;

// group attributes:
	  :data_provider = "/home/huanwu/summa/fork/summa/setup_tools/input/" ;
	  :data_reference = "/home/huanwu/summa/fork/summa/setup_tools/output/" ;

data:

   HRUarea = 32700, 32700, 32700, 32700, 32700 ;

   latitude = 43.2, 43.2, 43.2, 43.2, 43.2 ;

   longitude = 243.2, 243.2, 243.2, 243.2, 243.2 ;

   elevation = 2097, 2097, 2097, 2097, 2097 ;

   tan_slope = 0.20826, 0.20826, 0.20826, 0.20826, 0.20826 ;

   contourLength = 180.83141, 180.83141, 180.83141, 180.83141, 180.83141 ;

   mHeight = 19.25, 19.25, 19.25, 19.25, 19.25 ;

  } // group hru_attributes
}
